module OIP_palette (
	input logic [7:0] index,
	output logic [3:0] red, green, blue
);

localparam [0:255][11:0] palette = {
	{4'hE, 4'hE, 4'hE},
	{4'hD, 4'hD, 4'hD},
	{4'hF, 4'hF, 4'hF},
	{4'hB, 4'hB, 4'hB},
	{4'hB, 4'hB, 4'hB},
	{4'hD, 4'hD, 4'hD},
	{4'h9, 4'h9, 4'h9},
	{4'hF, 4'hF, 4'hF},
	{4'hC, 4'hC, 4'hC},
	{4'hE, 4'hE, 4'hE},
	{4'hD, 4'hD, 4'hD},
	{4'hA, 4'hA, 4'hA},
	{4'hC, 4'hC, 4'hC},
	{4'hE, 4'hE, 4'hE},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hE, 4'hE, 4'hE},
	{4'hD, 4'hD, 4'hD},
	{4'hC, 4'hC, 4'hC},
	{4'h9, 4'h9, 4'h9},
	{4'hA, 4'hA, 4'hA},
	{4'hD, 4'hD, 4'hD},
	{4'hD, 4'hD, 4'hD},
	{4'hB, 4'hB, 4'hB},
	{4'hF, 4'hF, 4'hF},
	{4'hB, 4'hB, 4'hB},
	{4'hC, 4'hC, 4'hC},
	{4'hF, 4'hF, 4'hF},
	{4'hE, 4'hE, 4'hE},
	{4'hE, 4'hE, 4'hE},
	{4'hF, 4'hF, 4'hF},
	{4'hA, 4'hA, 4'hA},
	{4'hF, 4'hF, 4'hF},
	{4'hA, 4'hA, 4'hA},
	{4'hE, 4'hE, 4'hE},
	{4'h9, 4'h9, 4'h9},
	{4'hF, 4'hF, 4'hF},
	{4'hD, 4'hD, 4'hD},
	{4'hC, 4'hC, 4'hC},
	{4'hC, 4'hC, 4'hC},
	{4'h9, 4'h9, 4'h9},
	{4'hE, 4'hE, 4'hE},
	{4'hD, 4'hD, 4'hD},
	{4'hE, 4'hE, 4'hE},
	{4'hA, 4'hA, 4'hA},
	{4'hD, 4'hD, 4'hD},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hD, 4'hD, 4'hD},
	{4'hF, 4'hF, 4'hF},
	{4'hE, 4'hE, 4'hE},
	{4'hD, 4'hD, 4'hD},
	{4'hC, 4'hC, 4'hC},
	{4'hB, 4'hB, 4'hB},
	{4'hA, 4'hA, 4'hA},
	{4'hB, 4'hB, 4'hB},
	{4'hD, 4'hD, 4'hD},
	{4'hD, 4'hD, 4'hD},
	{4'h9, 4'h9, 4'h9},
	{4'hB, 4'hB, 4'hB},
	{4'hE, 4'hE, 4'hE},
	{4'hE, 4'hE, 4'hE},
	{4'hD, 4'hD, 4'hD},
	{4'hF, 4'hF, 4'hF},
	{4'hC, 4'hC, 4'hC},
	{4'hF, 4'hF, 4'hF},
	{4'hE, 4'hE, 4'hE},
	{4'hB, 4'hB, 4'hB},
	{4'hC, 4'hC, 4'hC},
	{4'hF, 4'hF, 4'hF},
	{4'hC, 4'hC, 4'hC},
	{4'hC, 4'hC, 4'hC},
	{4'hB, 4'hB, 4'hB},
	{4'hF, 4'hF, 4'hF},
	{4'hC, 4'hC, 4'hC},
	{4'hE, 4'hE, 4'hE},
	{4'hD, 4'hD, 4'hD},
	{4'hC, 4'hC, 4'hC},
	{4'hE, 4'hE, 4'hE},
	{4'hB, 4'hB, 4'hB},
	{4'hE, 4'hE, 4'hE},
	{4'hC, 4'hC, 4'hC},
	{4'hB, 4'hB, 4'hB},
	{4'hC, 4'hC, 4'hC},
	{4'hA, 4'hA, 4'hA},
	{4'hD, 4'hD, 4'hD},
	{4'hC, 4'hC, 4'hC},
	{4'hB, 4'hB, 4'hB},
	{4'h9, 4'h9, 4'h9},
	{4'hB, 4'hB, 4'hB},
	{4'hC, 4'hC, 4'hC},
	{4'hA, 4'hA, 4'hA},
	{4'hB, 4'hB, 4'hB},
	{4'hA, 4'hA, 4'hA},
	{4'hA, 4'hA, 4'hA},
	{4'hA, 4'hA, 4'hA},
	{4'hB, 4'hB, 4'hB},
	{4'h9, 4'h9, 4'h9},
	{4'hA, 4'hA, 4'hA},
	{4'h9, 4'h9, 4'h9},
	{4'hA, 4'hA, 4'hA},
	{4'hA, 4'hA, 4'hA},
	{4'hA, 4'hA, 4'hA},
	{4'hA, 4'hA, 4'hA},
	{4'h9, 4'h9, 4'h9},
	{4'hB, 4'hB, 4'hB},
	{4'h9, 4'h9, 4'h9},
	{4'h9, 4'h9, 4'h9},
	{4'h8, 4'h8, 4'h8},
	{4'hB, 4'hB, 4'hB},
	{4'hC, 4'hC, 4'hC},
	{4'hB, 4'hB, 4'hA},
	{4'hE, 4'hE, 4'hD},
	{4'hF, 4'hF, 4'hF},
	{4'hB, 4'hB, 4'hB},
	{4'hD, 4'hD, 4'hD},
	{4'h9, 4'h9, 4'h9},
	{4'hC, 4'hC, 4'hC},
	{4'hB, 4'hB, 4'hB},
	{4'h9, 4'h9, 4'h9},
	{4'h9, 4'h9, 4'h9},
	{4'hC, 4'hC, 4'hC},
	{4'hC, 4'hC, 4'hC},
	{4'hB, 4'hB, 4'hB},
	{4'hD, 4'hD, 4'hD},
	{4'hF, 4'hF, 4'hF},
	{4'hC, 4'hC, 4'hC},
	{4'hC, 4'hC, 4'hC},
	{4'hE, 4'hE, 4'hE},
	{4'hB, 4'hB, 4'hB},
	{4'hC, 4'hC, 4'hC},
	{4'h9, 4'h9, 4'h9},
	{4'hC, 4'hC, 4'hC},
	{4'hF, 4'hF, 4'hF},
	{4'hC, 4'hC, 4'hC},
	{4'hC, 4'hC, 4'hC},
	{4'hE, 4'hE, 4'hE},
	{4'hC, 4'hC, 4'hC},
	{4'hF, 4'hF, 4'hF},
	{4'hD, 4'hD, 4'hD},
	{4'hB, 4'hB, 4'hB},
	{4'hC, 4'hC, 4'hC},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF},
	{4'hF, 4'hF, 4'hF}
};

assign {red, green, blue} = palette[index];

endmodule
